library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.aes_pkg.all;

package aes_record_pkg is


	

end package aes_record_pkg;

package body aes_record_pkg is

end package body aes_record_pkg;
