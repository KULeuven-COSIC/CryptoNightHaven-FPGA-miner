`timescale 1 ps / 1 ps

module cryptonight(
  input  wire             ap_clk               ,          
  input  wire             ap_rst_n             ,
  output wire             interrupt            ,
  output wire     [63:0]  m00_axi_araddr       ,
  output wire     [1:0]   m00_axi_arburst      ,
  output wire     [3:0]   m00_axi_arcache      ,
  output wire     [7:0]   m00_axi_arlen        ,
  output wire     [0:0]   m00_axi_arlock       ,
  output wire     [2:0]   m00_axi_arprot       ,
  output wire     [3:0]   m00_axi_arqos        ,
  input  wire             m00_axi_arready      ,
  output wire     [2:0]   m00_axi_arsize       ,
  output wire             m00_axi_arvalid      ,
  output wire     [63:0]  m00_axi_awaddr       ,
  output wire     [1:0]   m00_axi_awburst      ,
  output wire     [3:0]   m00_axi_awcache      ,
  output wire     [7:0]   m00_axi_awlen        ,
  output wire     [0:0]   m00_axi_awlock       ,
  output wire     [2:0]   m00_axi_awprot       ,
  output wire     [3:0]   m00_axi_awqos        ,
  input  wire             m00_axi_awready      ,
  output wire     [2:0]   m00_axi_awsize       ,
  output wire             m00_axi_awvalid      ,
  output wire             m00_axi_bready       ,
  input  wire     [1:0]   m00_axi_bresp        ,
  input  wire             m00_axi_bvalid       ,
  input  wire     [127:0] m00_axi_rdata        ,
  input  wire             m00_axi_rlast        ,
  output wire             m00_axi_rready       ,
  input  wire     [1:0]   m00_axi_rresp        ,
  input  wire             m00_axi_rvalid       ,
  output wire     [127:0] m00_axi_wdata        ,
  output wire             m00_axi_wlast        ,
  input  wire             m00_axi_wready       ,
  output wire     [15:0]  m00_axi_wstrb        ,
  output wire             m00_axi_wvalid       ,
  input  wire     [11:0]  s_axi_control_araddr ,
  output wire             s_axi_control_arready,
  input  wire             s_axi_control_arvalid,
  input  wire     [11:0]  s_axi_control_awaddr ,
  output wire             s_axi_control_awready,
  input  wire             s_axi_control_awvalid,
  input  wire             s_axi_control_bready ,
  output wire     [1:0]   s_axi_control_bresp  ,
  output wire             s_axi_control_bvalid ,
  output wire     [31:0]  s_axi_control_rdata  ,
  input  wire             s_axi_control_rready ,
  output wire     [1:0]   s_axi_control_rresp  ,
  output wire             s_axi_control_rvalid ,
  input  wire     [31:0]  s_axi_control_wdata  ,
  output wire             s_axi_control_wready ,
  input  wire     [3:0]   s_axi_control_wstrb  ,
  input  wire             s_axi_control_wvalid 
  );

  cryptonight_bd inst_cryptonight_bd (.*);

endmodule